module test;
    initial begin
        $display("Verilog OK and ready.");
        $finish;
    end
endmodule